module qb(x1,x2,x3,x4,x5,f);
	input x1,x2,x3,x4,x5;
	output f;
	
