module encoder16to4(a,f);
	input [15:0] a;
	output reg [4:0] f;
	integer i;
	always @(a)
	begin
		for(i=0;i<16;i=i+1)
		begin
			
	end
endmodule
